entity somador8bits is 
end entity;
